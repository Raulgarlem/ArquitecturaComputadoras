contador12_inst : contador12 PORT MAP (
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		sclr	 => sclr_sig,
		sload	 => sload_sig,
		q	 => q_sig
	);
